module main (
	input A,
	output Z);

	assign Z =A;
endmodule
