module main ();

endmodule
